module branch_controller (
  input [31:0] inst,
  input cmpin,
  input pc,
  output addr_out,

);
